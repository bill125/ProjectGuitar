library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package definitions is
	subtype StringStatus is integer range 0 to 88;
	type GuitarStatus is array (0 to 5) of StringStatus;
end package	definitions;