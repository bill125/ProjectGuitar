entity Velocity is
  port (
	seg0, seg1 : in std_logic_vector(6 downto 0);
	vel : array (0 to 5) of integer
    );
end entity Velocity;

architecture beh of Velocity is
begin
  
end
